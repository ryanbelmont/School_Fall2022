parameter  LW = 6'b100011 ; 
parameter SW = 6'b101011 ;
parameter no_op = 32'b0000000_0000000_0000000_0000000 ;
parameter ALUop = 6'b0 ;
parameter CDEC = 6'b101111 ;
parameter IJMP=6'b110000 ;

string filename="/home/ryan/Documents/school/Fall2022/EE4363/EE4363_lab2/handout/specific_tests/IJMP/4/regs.dat";
string filename1="/home/ryan/Documents/school/Fall2022/EE4363/EE4363_lab2/handout/specific_tests/IJMP/4/dmem.dat";
string filename2="/home/ryan/Documents/school/Fall2022/EE4363/EE4363_lab2/handout/specific_tests/IJMP/4/imem.dat";
string filename3="/home/ryan/Documents/school/Fall2022/EE4363/EE4363_lab2/handout/specific_tests/IJMP/4/mem_result.dat";
string filename4="/home/ryan/Documents/school/Fall2022/EE4363/EE4363_lab2/handout/specific_tests/IJMP/4/regs_result.dat";

