parameter  LW = 6'b100011 ; 
parameter SW = 6'b101011 ;
parameter no_op = 32'b0000000_0000000_0000000_0000000 ;
parameter ALUop = 6'b0 ;
parameter CDEC = 6'b101111 ;
parameter IJMP=6'b110000 ;

string filename="regs.dat";
string filename1="dmem.dat";
string filename2="imem.dat";
string filename3="mem_result.dat";
string filename4="regs_result.dat";
