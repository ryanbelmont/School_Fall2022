`timescale 1ns / 1ps


module comparator_1b(A, B, less_or_eq);
    input A, B;
    output less_or_eq;
    
endmodule
