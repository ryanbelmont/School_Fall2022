`timescale 1ns / 1ps


module mux4to1(out, a, b, c, d, s0, s1);
    input a, b, c, d, s0, s1;
    output out;

endmodule
